module oauth1

pub fn generate_oauth1_header() string {
	return ""
}