module oauth1

pub struct Config {
pub mut:
	consumer_key string
	consumer_secret string
	call_back_url string
}